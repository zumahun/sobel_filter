module hdmi_mod(

);


endmodule