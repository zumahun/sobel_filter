module cam_ctrl(
    input sys_clk_i,
    input sys_rst_i,

    output xvclk_o,
    output sio_c_o,
    inout sio_d_io,

    output cam_rst_o,
    output cam_pwd_o
);


endmodule